module instruction_fetch
(input clk,
    
);

endmodule