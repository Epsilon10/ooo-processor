module instruction_buffer
(input clk,
input valid_0, input [3:0] opcode_0, input [3:0] r_a_0, input [3:0] r_b_0, input [3:0] rt_0,
input valid_1, input [3:0] opcode_1, input [3:0] r_a_1, input [3:0] r_b_1, input [3:0] rt_1,
input valid_2, input [3:0] opcode_2, input [3:0] r_a_2, input [3:0] r_b_2, input [3:0] rt_2,
input valid_3, input [3:0] opcode_3, input [3:0] r_a_3, input [3:0] r_b_3, input [3:0] rt_3,
);

endmodule